library ieee;
use ieee.std_logic_1164.all;

entity adder is
    port (a: in std_logic_vector (3 downto 0);
          in2 : in std_logic_vector (3 downto 0);
          sum : out std_logic_vector(3 downto 0));
end adder;

architecture sum of adder is


end sum;
